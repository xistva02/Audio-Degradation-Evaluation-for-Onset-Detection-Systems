BZh91AY&SYI�j$ �_�Py����߰����`�  ��    2dɈ��	�����q�&LF& L�&@F ���2b10d�2 h�00O�H         �zM24d�4F&#F�2 �$@A4�2i� �5	�4P&&�l��$��&$�p����)J]!�"�?W��>�U$UQQ(X��rJª��0D�%H?�C5!�X��:F�=:�*�]�N�&�v�\�IXޫ#Scői�N�j�T�UUJb��u���
M�z�3f��.�~	�zc���ʥR�^'������n����Y�ɪ�cư�)9�u�T������ra�}2����\#�8�2���ɕg���I:$`�v���{�K����>���qOҪ�N��5"��UJ���IIE(�Xg"q�o;�';��Ɋ�Ŋ���͊^�f��_�t.ŤC�z���(�+�S�I�سyQ��Sj��UJ��Ir��k�4d��b�L����B�6L5Yf�mQ�m-�X63b��&2��kk��&<��F�G1���oS�Y0f�u�'�t�;�%RR��   1�cI�+I1w=-A�RR��c,S�L�Q�=�x.���꾌ZT��M
eThY��R�Y/{)B���/V^ԥ�{�K���V�ѵ�cr��b�,R5�o��UUN��(�6V�E���N���S�lR�	� 0���> uh��$�̳���iy����Cbj�K�v=�#݄h��x�#c�'�F�C�y���	��?I�O|��%��#bv�z��s������,>	g��u攛����G���X0>j)q�)cd�6$Y>F�UT.�R>�M,����0(��-�9�\��X�o.���͡��:��RN���iLB�s��T��H����KYw��sCP����>�mK!��c�'Y��)53z&�s�"�N�ނsM��ԣ`O�1��{d?���X��w)'�^G'j<f'����E9.QL�X6�$��zx�C���0:ʆ�A;����5�<�1�F�:�Vr~�$S�l_#�(�L��mN4�N�>��"�s�G��GYK�'!�܅��9��$�/!�!�b�0sҢ�K�E7�XKAD��:^$���4`�J,�T�kG%̢L�i#��a�EH���f�`Q��C��K#�9���k �]H�=# ~/#��������}Gy��O�4<��g<�������t����:��19*�����O4]#R�%���*T�i���G\~���3'[sQ�l�ԑ�7
c#�&*��IhS��,�E��N���)J\�;$b�ӗf֥Z���"�,v�EɈ�/��X��֣S����i�#��A���]I�bM瓉���dMZ��,dd.1�X~��07�sʉ���h^7�:�*]��:���oY�YLh����thOw�gINՖ���P6S���]��BA'ݨ�