BZh91AY&SY��c= �߀Py����߰����`
_<��:g@ M�yT*I(P��z�� 4ѐ�d=@���4�Q4�=   �  ��b�LFCC �#	5$�B�12hɐhh�C�(�hDbb5G�z�az�OH���i6��?SQ����4�� �@�˨F'�t�Z-��ݫ��O[,�h��I�>���,-lI�1�	� �Q!�^R�U��.�^FH��$b�I2!0`n��yjT�o��� w�x�O��r��ٖP��!�0�a�Z��m}XL�Q���5�L��x��7s�.�nG��x��ܜ�&
S�@�V�qޫ5Dl8(`�}sR��]�Nj"!`J�xkn�?��y. ���E��Q���|�ٴe�G&���#���6M��M�Kk2 �p���[�VϹAd6���	�7�x��(Ѕ5�A�:C��v���G���c����ݫ�ǀw'��#�@jw{��gFhZ��C��T�KQ�������plڤ��V���9:�昩8,<����"�v0f((؁�Μ�n1`6��4@a���do͖��Å�g�=t��@�i�B�=?�$��߅��WYd&�j`uXu�@��Pً�S� ML��`[�ꥵ.[W%U�M�0-�1�I3��<!���j\����?0v 7z`H몇Oǐ�����P.��D���	��$n�`�CW�ӊ��պ�8�R�Ƈ�0YܻUhi�j|� �A�I���p1
3��Z)q�pc���=(�i�u}�p
ͧX�7p�h�k�d��s3-��j!�%h"1k�pi��.�������Q��p�t�eF�����3\���R�n�pp��J"�B9ɲ��)kQ�{MH��r2����g����o�`1N��=���-q�řy�37)�"��ppK�	�_u�r��Ы�:�yXx.��Bav#﷎qO�<�H�F.�UUUUUB! (������)K�́����X(56���ƭ�LSh����K�B�F#b �IG],�)���SH�k%�P@�]k]IR֠-IR�P,�����4CF̺�C6A��s�=Zj��J�� E�d��Tҏ���:���V����F �&:�"� "�(	����h;Z�N<P��|8>�{��.O0����p���
��ߵ��C���HU���(��B�����=>@�t��%�G G�p,,�Qw�]���t#�b5/4b��y#1ϲ����</j!���E=�� `��x?&y�=�!G	'�P*�1ML%�9�!�m�Ys�n�0�]
:���[žy��k���;�ɳ,4v�e
#�ܛ?[/[G6�XEe�!����#G��!��.��Qԅ�wV��kn�j��!̵^he�m�,��#m�<c����l�ż�W u�c���`h����s�/��w�nx�`�K�2]wv1j�����jrC�>�g�K.k"��(K��n;ֈt��`ty��tg5�m�X��'�zP �kCqB$bW�;A��pJv!���}�`��̸���v�,��5q���c�W{� �(s(�4B���Z���-��a�+1��B�ͽn�	2]���j�9���K�.cQ��,����h� ]P�a�,�P�&�7*֬��j�Pe'��<�r��W�-`�n�|r�m��e����.۲䆞�k�:������PWS�2�����zی>�x0�y����=������im��{уo���^� *���}C���Hf� ��]@�d9������@�db�d=MYz��(�w�]Ɂ�ɨ�:��nb��,A��0Ψ `��r�\#�o�3a�,=�twۋ�s�#D,ё�7�s�ͻ�:990��n�j*���@0��� ?�%܇��h<ʇ�`���������A��ha]ýcw?.֏H��� �`@,�������H�
<Lg�